import fpnew_pkg::*; 

package expu_pkg;
    typedef enum int unsigned { BEFORE, AFTER, AROUND } regs_config_t;
endpackage