import fpnew_pkg::*;

package sfm_pkg;
    typedef enum int unsigned { BEFORE, AFTER, AROUND } regs_config_t;
    typedef enum int unsigned { MIN, MAX }              min_max_mode_t;

    function sfm_to_cvfpu(sfm_pkg::regs_config_t arg);
        fpnew_pkg::pipe_config_t res;

        unique case (arg)
            sfm_pkg::BEFORE :   res = fpnew_pkg::BEFORE;
            sfm_pkg::AFTER  :   res = fpnew_pkg::AFTER;
            sfm_pkg::AROUND :   res = fpnew_pkg::DISTRIBUTED;
        endcase

        return res;
    endfunction
endpackage